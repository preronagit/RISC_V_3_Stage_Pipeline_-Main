module tb();

    reg clk=0, rst;
    Pipeline_top pipeline (.clk(clk), .rst(rst));
    always begin
        clk = ~clk;
        #50;
    end

    initial begin
        rst <= 1'b0;
        #200;
        rst <= 1'b1;
        #1000;
        $finish;    
    end

    initial begin
        $dumpfile("pipeline_3_stage.vcd");
        $dumpvars(0);
    end

   
endmodule